// Global variables
int nop;
int nop_out;
int error;